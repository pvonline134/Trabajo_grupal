module binary_to_7segm (

    input logic [3:0] binary,
    output logic [6:0] segments,

);
    
endmodule
    
    

